`timescale 1ns / 1ps

module npc(
    input [31:0] PC,
	 input [31:0] RA,
    input [25:0] Imm,
    input [1:0] NPCOp,
    output [31:0] PC4,
    output [31:0] NPC
    );

    //PC4
    assign PC4 = PC + 4;

    //ALUOp determines NPC
    assign NPC = (NPCOp == 2'b00) ? PC + 4 :                               	   // sequense execution
                 (NPCOp == 2'b01) ? PC + 4 + {{14{Imm[15]}}, Imm[15:0], 2'b0} :  // conditional branch (PC + 4 + offset), sign extend!!!
                 (NPCOp == 2'b10) ? {PC[31:28], Imm, 2'b0} :                     // unconditional jump
                 RA;           

endmodule
